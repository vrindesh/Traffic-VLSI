//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/03/2024 12:06:23 AM
// Design Name: 
// Module Name: final
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module final(input clk,output [0:2]r,[0:2]g,[0:2]y );
//reg [0:4]Q;
//reg [0:31]s;
//always@(clk)
//begin
//counterc1 (clk,Q[0],Q[1],Q[2],Q[3] );
//demuxd1  (
//end
//endmodule
